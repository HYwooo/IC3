
module KeyToDigits (
    
);
    
endmodule